module four_bit_adder(a,b,s,c);
input [3:0]a;
input [3:0]b;

output [3:0]s;
output [3:0]c;

assign s = a^b;
assign c = a&b;

endmodule 